



// class sequncer

class destin_seqr extends uvm_sequencer#(destin_xtn);

// factory registration

         `uvm_component_utils(destin_seqr)

// function new constructor

		 function new(string name = "destin_seqr",uvm_component parent);
		 
				super.new(name,parent);
		 
		 endfunction







endclass