

// source xtn

class source_xtn extends uvm_sequence_item;

// factory registration

		`uvm_object_utils(source_xtn)

	  		

// function new

		function new(string name = "source_xtn");
		
				super.new(name);
		
		endfunction


endclass