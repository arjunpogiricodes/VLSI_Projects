



// class sequncer

class source_seqr extends uvm_sequencer#(source_xtn);

// factory registration

         `uvm_component_utils(source_seqr)

// function new constructor

		 function new(string name = "source_seqr",uvm_component parent);
		 
				super.new(name,parent);
		 
		 endfunction







endclass