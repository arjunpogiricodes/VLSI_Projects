

// source xtn

class destin_xtn extends uvm_sequence_item;

// factory registration

		`uvm_object_utils(destin_xtn)

// function new

		function new(string name = "destin_xtn");
		
				super.new(name);
		
		endfunction


endclass