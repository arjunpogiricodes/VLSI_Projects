

// --------- ahb to apb packages ------------------//

package ahbtoapb_pkg;

       import uvm_pkg::*;
       `include "uvm_macros.svh"
       `include "definitions.v"

       `include "ahb_config.sv"
       `include "apb_config.sv"

       `include "tb_env_config.sv"

       `include "apb_xtn.sv"
       `include "ahb_xtn.sv"

       `include "ahb_drvier.sv"
       `include "ahb_monitor.sv"
       `include "ahb_seqr.sv"
       `include "ahb_seq.sv"
       `include "ahb_agent.sv"
       `include "ahb_agent_top.sv"

       `include "apb_driver.sv"
       `include "apb_monitor.sv"
       `include "apb_seqr.sv"
       `include "apb_seq.sv"
       `include "apb_agent.sv"
       `include "apb_agent_top.sv"
       `include "virtual_seqr.sv"
       `include "virtual_seq.sv" 
       `include "tb_scoreboard.sv"
       `include "tb_env.sv"
       `include "base_test.sv"

endpackage
